/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
///Q=======================================================
//  MODULE Definition
//=======================================================
module CC_MUX3 #(parameter MUX3_SELECTWIDTH=2,parameter MUX3_NADAWIDTH=8, parameter MUX3_UBICACIONWIDTH=8)(
//////////// OUTPUTS //////////
	CC_POSICION_Out,
//////////// INPUTS //////////
	CC_MUX3_select_InBUS,
	CC_MUX3_NADA_InBUS,
	CC_MUX3_UBICACION_InBUS
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output	reg CC_POSICION_Out;
input 	[MUX3_SELECTWIDTH-1:0] CC_MUX3_select_InBUS;
input 	[MUX3_NADAWIDTH-1:0] CC_MUX3_NADA_InBUS;
input 	[MUX3_UBICACIONWIDTH-1:0] CC_MUX3_UBICACION_InBUS;
//=======================================================Q/
///A=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
always @(CC_MUX3_NADA_InBUS or CC_MUX3_UBICACION_InBUS or CC_MUX3_select_InBUS)
begin
   if( CC_MUX3_select_InBUS == 0)
      CC_POSICION_Out = CC_MUX3_UBICACION_InBUS;
   else if( CC_MUX3_select_InBUS == 1)
      CC_POSICION_Out = CC_MUX3_NADA_InBUS;
end

endmodule