/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
///Q=======================================================
//  MODULE Definition
//=======================================================
module CC_MUX12 #(parameter MUX12_SELECTWIDTH=2,parameter MUX12_NADAWIDTH=8, parameter MUX12_RANDOM1WIDTH=8, parameter MUX12_RANDOM2WIDTH=8, parameter MUX12_RANDOM3WIDTH=8 )(
//////////// OUTPUTS //////////
	CC_SALIDARANDOMS_Out,
//////////// INPUTS //////////
	CC_MUX12_select_InBUS,
	CC_MUX12_NADA_InBUS,
	CC_MUX12_RANDOM1_InBUS,
	CC_MUX12_RANDOM2_InBUS,
	CC_MUX12_RANDOM3_InBUS
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output	reg [MUX12_NADAWIDTH-1:0]CC_SALIDARANDOMS_Out;
input 	[MUX12_SELECTWIDTH-1:0] CC_MUX12_select_InBUS;
input 	[MUX12_NADAWIDTH-1:0] CC_MUX12_NADA_InBUS;
input 	[MUX12_RANDOM1WIDTH-1:0] CC_MUX12_RANDOM1_InBUS;
input 	[MUX12_RANDOM2WIDTH-1:0] CC_MUX12_RANDOM2_InBUS;
input 	[MUX12_RANDOM3WIDTH-1:0] CC_MUX12_RANDOM3_InBUS;
//=======================================================Q/
///A=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
always @(*)
begin
   if( CC_MUX12_select_InBUS == 0)
      CC_SALIDARANDOMS_Out = CC_MUX12_NADA_InBUS;
   else if( CC_MUX12_select_InBUS == 1)
      CC_SALIDARANDOMS_Out = CC_MUX12_RANDOM1_InBUS;
   else if( CC_MUX12_select_InBUS == 2)
      CC_SALIDARANDOMS_Out = CC_MUX12_RANDOM2_InBUS;
   else //if( CC_MUX12_select_InBUS == 3)
      CC_SALIDARANDOMS_Out = CC_MUX12_RANDOM3_InBUS;
end

endmodule