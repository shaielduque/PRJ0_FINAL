/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
///Q=======================================================
//  MODULE Definition
//=======================================================
module CC_MUX11 #(parameter MUX11_SELECTWIDTH=1,parameter MUX11_NADAWIDTH=8, parameter MUX11_TRANSIWIDTH=8)(
//////////// OUTPUTS //////////
	CC_TRANSI3_Out,
//////////// INPUTS //////////
	CC_MUX11_select_InBUS,
	CC_MUX11_NADA_InBUS,
	CC_MUX11_TRANSI_InBUS
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
output	reg CC_TRANSI3_Out;
input 	[MUX11_SELECTWIDTH-1:0] CC_MUX11_select_InBUS;
input 	[MUX11_NADAWIDTH-1:0] CC_MUX11_NADA_InBUS;
input 	[MUX11_TRANSIWIDTH-1:0] CC_MUX11_TRANSI_InBUS;
//=======================================================Q/
///A=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
always @(CC_MUX11_NADA_InBUS or CC_MUX11_TRANSI_InBUS or CC_MUX11_select_InBUS)
begin
   if( CC_MUX11_select_InBUS == 0)
      CC_TRANSI3_Out = CC_MUX11_TRANSI_InBUS;
   else if( CC_MUX11_select_InBUS == 1)
      CC_TRANSI3_Out = CC_MUX11_TRANSI_InBUS;
end

endmodule